// Copyright(C) 2019-2020 Lars Pontoppidan. All rights reserved.
// Use of this source code is governed by an MIT license file distributed with this software package
module java

pub const (
	keywords = [
		'abstract',
		'assert',
		'boolean',
		'break',
		'byte',
		'case',
		'catch',
		'char',
		'class',
		'const',
		'continue',
		'default',
		'do',
		'double',
		'else',
		'enum',
		'extends',
		'final',
		'finally',
		'float',
		'for',
		'goto',
		'if',
		'implements',
		'import',
		'instanceof',
		'int',
		'interface',
		'long',
		'native',
		'new',
		'package',
		'private',
		'protected',
		'public',
		'return',
		'short',
		'static',
		'strict',
		'super',
		'switch',
		'synchronized',
		'this',
		'throw',
		'throws',
		'transient',
		'try',
		'void',
		'volatile',
		'while',
	]
)
