// Copyright(C) 2019-2024 Lars Pontoppidan. All rights reserved.
// Use of this source code is governed by an MIT license file distributed with this software package
// This module handles everything related to user commands.
module user

import os
import compress.szip
import vab.paths
import vab.vxt
import net.http

const valid_sources = ['github']
pub const command_prefix = 'vab'

@[params]
pub struct InstallOptions {
pub:
	input     []string
	verbosity int
}

pub struct Command {
pub:
	id     string
	source string
	unit   string
	exe    string
}

// verbose prints `msg` to STDOUT if `InstallOptions.verbosity` level is >= `verbosity_level`.
pub fn (io &InstallOptions) verbose(verbosity_level int, msg string) {
	if io.verbosity >= verbosity_level {
		println(msg)
	}
}

// run_command runs a user installed command if found in `args`.
// If the command is found this function will call `exit()` with the result
// returned by the executed command.
pub fn run_command(args []string) {
	// Indentify user installed commands
	user_commands := commands()
	for _, user_command in user_commands {
		if user_command.id.trim_left('${command_prefix}-') in args {
			// First encountered known sub-command is executed on the spot.
			exit(launch_command(args[args.index(user_command.id.trim_left('${command_prefix}-'))..]))
		}
	}
}

fn launch_command(args []string) int {
	mut cmd := args[0]
	user_commands := commands()
	if command := user_commands['${command_prefix}-' + cmd] {
		tool_args := args[1..].clone()
		tool_exe := command.exe
		if os.is_executable(tool_exe) {
			// os.setenv('VAB_EXE', os.join_path(exe_dir, exe_name), true)
			$if windows {
				exit(os.system('${os.quoted_path(tool_exe)} ${tool_args}'))
			} $else $if js {
				// no way to implement os.execvp in JS backend
				exit(os.system('${tool_exe} ${tool_args}'))
			} $else {
				os.execvp(tool_exe, tool_args) or { panic(err) }
			}
			exit(2)
		}
		exec := (tool_exe + ' ' + tool_args.join(' ')).trim_right(' ')
		eprintln(@MOD + '.' + @FN + ' failed executing "${exec}"')
		return 1
	}

	eprintln(@MOD + '.' + @FN + ' failed to identify "${args}"')
	return 1
}

// install_command retrieves, installs and registers external user commands
pub fn install_command(opt InstallOptions) ! {
	// `vab install cmd xyz/abc`
	if opt.input.len == 0 {
		return error('${@FN} requires input')
	}

	component := opt.input[0] // Only 1 argument needed for now

	if component.count(':') == 0 {
		// no source protocol detected, slap on default and try again...
		mod_opt := InstallOptions{
			...opt
			input: ['github:${component}']
		}
		return install_command(mod_opt)
	}

	source := component.all_before(':')
	if source !in valid_sources {
		return error('${@FN} unknown source `${source}`. Valid sources are ${valid_sources}')
	}
	unit := component.all_after(':')

	match source {
		'github' {
			return install_from_github(unit, opt.verbosity)
		}
		else {
			return error('${@FN} unknown source `${source}`. Valid sources are ${valid_sources}')
		}
	}
}

fn install_from_github(unit string, verbosity int) ! {
	if unit.count('/') != 1 {
		return error('${@MOD} ${@FN} `${unit}` should contain exactly one "/" character')
	}
	unit_parts := unit.split('/')

	// TODO: support @ notation for specific commits/branches?
	// mut at_part := unit.all_after('@')

	if !(valid_identifier(unit_parts[0]) && valid_identifier(unit_parts[1])) {
		return error('${@MOD} ${@FN} `${unit}` is not a valid identifier')
	}
	initial_dst := os.join_path(paths.cache(), 'user', 'commands', 'github', unit_parts[0]) // TODO: const these

	url := 'https://github.com/${unit}/archive/refs/heads/master.zip'
	tmp_downloads := os.join_path(paths.tmp_work(), 'user', 'downloads') // TODO: const these
	paths.ensure(tmp_downloads)!

	zip_file := os.join_path(tmp_downloads, 'github-${unit.replace('/', '-')}.zip')
	if !os.exists(zip_file) {
		if verbosity > 1 {
			println('Downloading `${unit}` from "${url}"...')
		}
		http.download_file(url, zip_file) or {
			return error('${@MOD} ${@FN} failed to download `${unit}`: ${err}')
		}
	}
	final_dst := os.join_path(initial_dst, unit_parts[1])
	// Install
	if verbosity > 1 {
		println('Installing `${unit}` to "${final_dst}"...')
	}
	paths.ensure(initial_dst)!

	unzip(zip_file, initial_dst)!
	unzipped_dst := os.join_path(initial_dst, '${unit_parts[1]}-master')
	if os.exists(final_dst) {
		os.rmdir_all(final_dst) or {}
	}
	os.mv(unzipped_dst, final_dst)!

	build_command(final_dst, verbosity)!
	record_install(unit_parts[1], 'github', unit)!
}

fn record_install(id string, source string, unit string) ! {
	path := os.join_path(paths.cache(), 'user') // TODO: const these
	paths.ensure(path)!
	installs_db := os.join_path(path, 'installed.txt') // TODO: const these
	installs_db_bak := os.join_path(path, 'installed.txt.bak') // TODO: const these
	if !os.exists(installs_db) {
		os.create(installs_db)!
	}
	mut installs := os.read_lines(installs_db)!

	mut found := false
	for install_line in installs {
		if install_line == '' || install_line.starts_with('#') {
			continue
		}
		split := install_line.split(';')
		if split.len > 0 {
			if split[0] == id {
				found = true
				break
			}
		}
	}
	if !found {
		installs << '${id};${source};${unit}'
		os.mv(installs_db, installs_db_bak, overwrite: true)!
		os.write_lines(installs_db, installs)!
	}
}

pub fn has(command string) bool {
	cmds := commands()
	return command in cmds.keys()
}

pub fn commands() map[string]Command {
	mut installed := map[string]Command{}
	path := os.join_path(paths.cache(), 'user') // TODO: const these
	installs_db := os.join_path(path, 'installed.txt') // TODO: const these
	if os.exists(installs_db) {
		installs := os.read_lines(installs_db) or { return installed }
		for install_line in installs {
			if install_line == '' || install_line.starts_with('#') {
				continue
			}
			split := install_line.split(';')
			if split.len > 2 {
				id := split[0]
				source := split[1] or { 'unknown' }
				unit := split[2] or { 'unknown/unknown' }
				unit_parts := unit.split('/')
				// TODO: support @ notation for specific commits/branches?
				// mut at_part := unit.all_after('@')
				final_dst := os.join_path(paths.cache(), 'user', 'commands', source, unit_parts[0],
					unit_parts[1]) // TODO: const these

				installed[id] = Command{
					id:     split[0]
					source: source
					unit:   unit
					exe:    os.join_path(final_dst, id)
				}
			}
		}
	}
	return installed
}

fn unzip(file string, dir string) ! {
	if !os.is_dir(dir) {
		os.mkdir_all(dir)!
	}
	szip.extract_zip_to_dir(file, dir)!
}

fn valid_identifier(s string) bool {
	if s.len == 0 {
		return false
	}
	for ch in s {
		if !(ch.is_letter() || ch.is_digit() || ch == `_` || ch == `-`) {
			return false
		}
	}
	return true
}

fn build_command(path string, verbosity int) ! {
	if !vxt.found() {
		return error('${@MOD} ${@FN} failed to locate a V compiler')
	}
	v_exe := vxt.vexe()
	v_cmd := [
		v_exe,
		path,
	]
	verbosity_print_cmd(v_cmd, verbosity)
	res := run(v_cmd)
	if res.exit_code != 0 {
		return error('${@MOD} ${@FN} "${v_cmd.join(' ')}" failed:\n${res.output}')
	}
}

// verbosity_print_cmd prints information about the `args` at certain `verbosity` levels.
fn verbosity_print_cmd(args []string, verbosity int) {
	if args.len > 0 && verbosity > 1 {
		cmd_short := args[0].all_after_last(os.path_separator)
		mut output := 'Running ${cmd_short} From: ${os.getwd()}'
		if verbosity > 2 {
			output += '\n' + args.join(' ')
		}
		println(output)
	}
}

fn run(args []string) os.Result {
	res := os.execute(args.join(' '))
	return res
}
